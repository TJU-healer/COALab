`include "defines.v"

module id_stage(
    input  wire                     cpu_rst_n,
    
    // ��ȡָ�׶λ�õ�PCֵ
    input  wire [`INST_ADDR_BUS]    id_pc_i,

    // ��ָ��洢��������ָ����?
    input  wire [`INST_BUS     ]    id_inst_i,

    // ��ͨ�üĴ����Ѷ��������� 
    input  wire [`REG_BUS      ]    rd1,
    input  wire [`REG_BUS      ]    rd2,

    //��ִ�н׶λ�õ�д���ź�?
    input wire                      exe2id_wreg,
    input wire [`REG_ADDR_BUS  ]    exe2id_wa,
    input wire [`REG_BUS       ]    exe2id_wd,

    //�ӷô�׶λ�õ�д����Ϣ
    input wire                      mem2id_wreg,
    input wire [`REG_ADDR_BUS  ]    mem2id_wa,
    input wire [`REG_BUS       ]    mem2id_wd,

    //��ִ�н׶κͷô�׶λش��Ĵ洢�����Ĵ�����ʹ���ź�?
    input wire                      exe2id_mreg,
    input wire                      mem2id_mreg,
      
    // ����ִ�н׶ε�������Ϣ
    output wire [`ALUTYPE_BUS  ]    id_alutype_o,
    output wire [`ALUOP_BUS    ]    id_aluop_o,
    output wire [`REG_ADDR_BUS ]    id_wa_o,
    output wire                     id_wreg_o,
    output wire                     id_whilo_o,   //дhilo�Ĵ���ʹ��
    output wire                     id_mreg_o,  

    // ����ִ�н׶ε�Դ������1��Դ������2
    output wire [`REG_BUS      ]    id_src1_o,
    output wire [`REG_BUS      ]    id_src2_o,
    output wire [`DATA_BUS     ]    id_din_o,
    output wire [`REG_BUS      ]    id_retaddr_o,
      
    // ������ͨ�üĴ����Ѷ˿ڵ�ʹ�ܺ͵�ַ
    output wire                     rreg1,
    output wire [`REG_ADDR_BUS ]    ra1,
    output wire                     rreg2,
    output wire [`REG_ADDR_BUS ]    ra2,
    
    output wire [ 1:0          ]    jtsel,
    output wire [`REG_BUS      ]    jump_addr_1,
    output wire [`REG_BUS      ]    jump_addr_2,
    output wire [`REG_BUS      ]    jump_addr_3,
    
    output wire                     stallreq_id,      //����׶η�������ͣ�����ź�?
    
    input  wire                     id_in_delay_i,    //��������׶ε�ָ�����ӳٲ�ָ��?
    input  wire                     flush_im,         //��մ�ָ��洢��������ָ��
    output wire [`REG_ADDR_BUS ]    cp0_addr,         //cp0�Ĵ����ĵ�ַ
    output wire [`INST_ADDR_BUS]    id_pc_o,          //��������׶ε�ָ���pcֵ
    output wire                     id_in_delay_o,    //��������׶ε�ָ�����ӳٲ�ָ��?
    output wire                     next_delay_o,     //��һ����������׶ε�ָ�����ӳٲ�ָ��?
    output wire [`EXC_CODE_BUS ]    id_exccode_o      //��������׶ε�ָ����쳣����
    );
    
    assign id_pc_o       = (cpu_rst_n == `RST_ENABLE) ? `PC_INIT : id_pc_i;
    assign id_in_delay_o = (cpu_rst_n == `RST_ENABLE) ? `FALSE_V : id_in_delay_i;
    
    // ����С��ģʽ��ָ֯����
    //�������ź�flush_im == 1����ȡ����ָ��Ϊ��ָ��
    wire [`INST_BUS] id_inst = (flush_im == `FLUSH) ? `ZERO_WORD : {id_inst_i[7:0], id_inst_i[15:8], id_inst_i[23:16], id_inst_i[31:24]};
    // wire [`INST_BUS] id_inst = (flush_im == `FLUSH) ? `ZERO_WORD : id_inst_i;

    // ��ȡָ�����и����ֶε���Ϣ
    wire [5 :0] op   = id_inst[31:26];
    wire [5 :0] func = id_inst[5 : 0];
    wire [4 :0] rd   = id_inst[15:11];
    wire [4 :0] rs   = id_inst[25:21];
    wire [4 :0] rt   = id_inst[20:16];
    wire [4 :0] sa   = id_inst[10: 6];
    wire [15:0] imm  = id_inst[15: 0]; 
    wire [25:0] instr_index = id_inst[25:0];

    /*-------------------- ��һ�������߼���ȷ����ǰ��Ҫ�����ָ��? --------------------*/
    wire inst_reg    = ~|op;
    wire inst_and    = inst_reg &  func[5] & ~func[4] & ~func[3] &  func[2] & ~func[1] & ~func[0];
    
    wire inst_subu   = inst_reg &  func[5] & ~func[4] & ~func[3] & ~func[2] &  func[1] &  func[0];
    wire inst_slt    = inst_reg &  func[5] & ~func[4] &  func[3] & ~func[2] &  func[1] & ~func[0];
    wire inst_add    = inst_reg &  func[5] & ~func[4] & ~func[3] & ~func[2] & ~func[1] & ~func[0];
    wire inst_mult   = inst_reg & ~func[5] &  func[4] &  func[3] & ~func[2] & ~func[1] & ~func[0];
    wire inst_mfhi   = inst_reg & ~func[5] &  func[4] & ~func[3] & ~func[2] & ~func[1] & ~func[0];
    wire inst_mflo   = inst_reg & ~func[5] &  func[4] & ~func[3] & ~func[2] &  func[1] & ~func[0];
    wire inst_sll    = inst_reg & ~func[5] & ~func[4] & ~func[3] & ~func[2] & ~func[1] & ~func[0];
    wire inst_ori    = ~op[5] & ~op[4] &  op[3] &  op[2] & ~op[1] &  op[0];
    wire inst_lui    = ~op[5] & ~op[4] &  op[3] &  op[2] &  op[1] &  op[0];
    wire inst_addiu  = ~op[5] & ~op[4] &  op[3] & ~op[2] & ~op[1] &  op[0];
    wire inst_sltiu  = ~op[5] & ~op[4] &  op[3] & ~op[2] &  op[1] &  op[0];
    wire inst_lb     =  op[5] & ~op[4] & ~op[3] & ~op[2] & ~op[1] & ~op[0];
    wire inst_lw     =  op[5] & ~op[4] & ~op[3] & ~op[2] &  op[1] &  op[0];
    wire inst_sb     =  op[5] & ~op[4] &  op[3] & ~op[2] & ~op[1] & ~op[0];
    wire inst_sw     =  op[5] & ~op[4] &  op[3] & ~op[2] &  op[1] &  op[0];
   
    wire inst_addu   = inst_reg &  func[5] & ~func[4] & ~func[3] & ~func[2] & ~func[1] &  func[0];
    wire inst_sub    = inst_reg &  func[5] & ~func[4] & ~func[3] & ~func[2] &  func[1] & ~func[0];
    wire inst_sltu   = inst_reg &  func[5] & ~func[4] &  func[3] & ~func[2] &  func[1] &  func[0];
    wire inst_or     = inst_reg &  func[5] & ~func[4] & ~func[3] &  func[2] & ~func[1] &  func[0];
    wire inst_nor    = inst_reg &  func[5] & ~func[4] & ~func[3] &  func[2] &  func[1] &  func[0];
    wire inst_xor    = inst_reg &  func[5] & ~func[4] & ~func[3] &  func[2] &  func[1] & ~func[0];
    wire inst_srl    = inst_reg & ~func[5] & ~func[4] & ~func[3] & ~func[2] &  func[1] & ~func[0];
    wire inst_sra    = inst_reg & ~func[5] & ~func[4] & ~func[3] & ~func[2] &  func[1] &  func[0];
    wire inst_sllv   = inst_reg & ~func[5] & ~func[4] & ~func[3] &  func[2] & ~func[1] & ~func[0];
    wire inst_srlv   = inst_reg & ~func[5] & ~func[4] & ~func[3] &  func[2] &  func[1] & ~func[0];
    wire inst_srav   = inst_reg & ~func[5] & ~func[4] & ~func[3] &  func[2] &  func[1] &  func[0];
    wire inst_multu  = inst_reg & ~func[5] &  func[4] &  func[3] & ~func[2] & ~func[1] &  func[0];
    wire inst_mthi   = inst_reg & ~func[5] &  func[4] & ~func[3] & ~func[2] & ~func[1] &  func[0];
    wire inst_mtlo   = inst_reg & ~func[5] &  func[4] & ~func[3] & ~func[2] &  func[1] &  func[0];
    wire inst_addi   = ~op[5] & ~op[4] &  op[3] & ~op[2] & ~op[1] & ~op[0];
    wire inst_slti   = ~op[5] & ~op[4] &  op[3] & ~op[2] &  op[1] & ~op[0];
    wire inst_andi   = ~op[5] & ~op[4] &  op[3] &  op[2] & ~op[1] & ~op[0];
    wire inst_xori   = ~op[5] & ~op[4] &  op[3] &  op[2] &  op[1] & ~op[0];
    wire inst_lbu    =  op[5] & ~op[4] & ~op[3] &  op[2] & ~op[1] & ~op[0];
    wire inst_lh     =  op[5] & ~op[4] & ~op[3] & ~op[2] & ~op[1] &  op[0];
    wire inst_lhu    =  op[5] & ~op[4] & ~op[3] &  op[2] & ~op[1] &  op[0];
    wire inst_sh     =  op[5] & ~op[4] &  op[3] & ~op[2] & ~op[1] &  op[0];
    
    wire inst_j      = ~op[5] & ~op[4] & ~op[3] & ~op[2] &  op[1] & ~op[0];
    wire inst_jal    = ~op[5] & ~op[4] & ~op[3] & ~op[2] &  op[1] &  op[0];
    wire inst_jr     = inst_reg & ~func[5] & ~func[4] &  func[3] & ~func[2] & ~func[1] & ~func[0];
    wire inst_beq    = ~op[5] & ~op[4] & ~op[3] &  op[2] & ~op[1] & ~op[0];
    wire inst_bne    = ~op[5] & ~op[4] & ~op[3] &  op[2] & ~op[1] &  op[0];
    
    wire inst_jalr   = inst_reg & ~func[5] & ~func[4] &  func[3] & ~func[2] & ~func[1] &  func[0];
    wire inst_bgez   = ~op[5]& ~op[4] & ~op[3] & ~op[2] & ~op[1] &  op[0] & ~id_inst[20] &  id_inst[16];
    wire inst_bgtz   = ~op[5]& ~op[4] & ~op[3] &  op[2] &  op[1] &  op[0];
    wire inst_blez   = ~op[5]& ~op[4] & ~op[3] &  op[2] &  op[1] & ~op[0];
    wire inst_bltz   = ~op[5]& ~op[4] & ~op[3] & ~op[2] & ~op[1] &  op[0] & ~id_inst[20] & ~id_inst[16];
    wire inst_bgezal = ~op[5]& ~op[4] & ~op[3] & ~op[2] & ~op[1] &  op[0] &  id_inst[20] &  id_inst[16];
    wire inst_bltzal = ~op[5]& ~op[4] & ~op[3] & ~op[2] & ~op[1] &  op[0] &  id_inst[20] & ~id_inst[16];
    
    wire inst_div    = inst_reg &~func[5]&  func[4] &  func[3] & ~func[2] &  func[1] & ~func[0];
    wire inst_divu   = inst_reg &~func[5]&  func[4] &  func[3] & ~func[2] &  func[1] &  func[0];    
    
    wire inst_syscall= inst_reg & ~func[5] & ~func[4] &  func[3] &  func[2] & ~func[1] & ~func[0];
    wire inst_eret   = ~op[5] &  op[4] & ~op[3] & ~op[2] & ~op[1] & ~op[0] & ~func[5]&  func[4] &  func[3] & ~func[2] & ~func[1] & ~func[0] ;
    wire inst_mfc0   = ~op[5] &  op[4] & ~op[3] & ~op[2] & ~op[1] & ~op[0] & ~id_inst[23];
    wire inst_mtc0   = ~op[5] &  op[4] & ~op[3] & ~op[2] & ~op[1] & ~op[0] &  id_inst[23];
    wire inst_break  = inst_reg & ~func[5] & ~func[4] &  func[3] &  func[2] & ~func[1] &  func[0];
    /*------------------------------------------------------------------------------*/

    /*-------------------- �ڶ��������߼������ɾ�������ź�? --------------------*/    
    wire rtsel  = (inst_addiu | inst_ori | inst_sltiu | inst_lui | inst_addi | inst_slti | inst_andi | inst_xori | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_sb | inst_sw | inst_sh | inst_mfc0);
    wire immsel = (inst_addiu | inst_ori | inst_sltiu | inst_lui | inst_addi | inst_slti | inst_andi | inst_xori | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_sb | inst_sw | inst_sh);
    wire sext   = (inst_addiu | inst_sltiu | inst_addi | inst_slti | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_sb | inst_sw | inst_sh);
    wire upper  = (inst_lui);
    wire jal    = (inst_jal | inst_bgezal | inst_bltzal);
    
    wire [`REG_BUS] imm_ext = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD :
                               (upper) ? imm << 16 :
                               (sext) ? { { 16 {imm[15]} }, imm} : {`ZERO_HWORD, imm};
                              
    wire [`REG_BUS] pc_next = id_pc_i + 4;
                               
    wire [1:0] fwrd1;
    wire [1:0] fwrd2;
    wire equ;
    
    // ��������alutype
    assign id_alutype_o[2] = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_sll | inst_srl | inst_sra | inst_sllv | inst_srlv | inst_srav | inst_j | inst_jal | inst_jr | inst_jalr | inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal | inst_syscall | inst_eret | inst_mtc0);
    assign id_alutype_o[1] = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_and | inst_ori | inst_lui | inst_andi | inst_nor | inst_or | inst_xor | inst_xori | inst_mfhi | inst_mflo | inst_syscall | inst_eret | inst_mfc0 | inst_mtc0 | inst_break);
    assign id_alutype_o[0] = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_add | inst_subu | inst_slt | inst_addiu | inst_sltiu | inst_addi | inst_addu | inst_sub | inst_slti | inst_sltu | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_sb | inst_sw | inst_sh | inst_mfhi | inst_mflo | inst_j | inst_jal | inst_jr | inst_jalr | inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal | inst_mfc0);

    // �ڲ�������aluop
    assign id_aluop_o[7]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (                                                                                                                                            inst_lb | inst_lw | inst_sb | inst_sw                                                                | inst_syscall | inst_eret | inst_mfc0 | inst_mtc0                                                                                                                                                                                                                                                                                               | inst_lh | inst_sh | inst_lbu | inst_lhu                        | inst_break); // 7
    assign id_aluop_o[6]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (                                                                                                                                                                                                                                                                                                      inst_addi | inst_addu | inst_sub                                                                                                                                        | inst_andi | inst_or | inst_xori                       | inst_sllv | inst_srlv | inst_srav                                                                                                      ); // 6                                                                                                                                                                                                                                                                                                                                     // 6
    assign id_aluop_o[5]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (                                  inst_slt                                                                        | inst_sltiu                                                    | inst_j | inst_jal | inst_jr | inst_beq | inst_bne                                                                                                  | inst_slti | inst_sltu              | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal                                                                                                                                                                                     | inst_jalr                        ); // 5
    assign id_aluop_o[4]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_add | inst_subu | inst_and |            inst_mult |                         inst_sll | inst_addiu | inst_ori                         | inst_lb | inst_lw | inst_sb | inst_sw                               | inst_beq | inst_bne | inst_div                                                                                                               | inst_multu | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal | inst_xor | inst_nor                                   | inst_srl | inst_sra                                                             | inst_lh | inst_sh | inst_lbu | inst_lhu             | inst_divu            ); // 4
    assign id_aluop_o[3]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_add | inst_subu | inst_and |                        inst_mfhi | inst_mflo |            inst_addiu | inst_ori                                             | inst_sb | inst_sw | inst_j | inst_jal | inst_jr                                                             | inst_mfc0 | inst_mtc0 | inst_addi | inst_addu | inst_sub | inst_slti | inst_sltu              | inst_bgez                                                                 | inst_xor | inst_nor | inst_andi | inst_or | inst_xori                                                           | inst_mthi | inst_mtlo           | inst_sh | inst_lbu | inst_lhu | inst_jalr                        ); // 3
    assign id_aluop_o[2]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (                       inst_and | inst_slt | inst_mult | inst_mfhi | inst_mflo |                         inst_ori | inst_sltiu | inst_lui                                         | inst_j | inst_jal | inst_jr                       | inst_div | inst_syscall | inst_eret | inst_mfc0 | inst_mtc0                                                            | inst_multu                                     | inst_bltz | inst_bgezal | inst_bltzal | inst_xor | inst_nor | inst_andi | inst_or | inst_xori                                                           | inst_mthi | inst_mtlo                                | inst_lhu | inst_jalr | inst_divu| inst_break); // 2
    assign id_aluop_o[1]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (           inst_subu |            inst_slt |                                                                        inst_sltiu                      | inst_lw           | inst_sw          | inst_jal                                 | inst_div | inst_syscall | inst_eret                                                 | inst_sub                                                  | inst_bgtz | inst_blez             | inst_bgezal | inst_bltzal | inst_xor | inst_nor                       | inst_xori | inst_srl | inst_sra             | inst_srlv | inst_srav | inst_mthi | inst_mtlo                     | inst_lbu            | inst_jalr | inst_divu            ); // 1
    assign id_aluop_o[0]   = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (           inst_subu |                                               inst_mflo | inst_sll | inst_addiu | inst_ori | inst_sltiu | inst_lui                                                             | inst_jr            | inst_bne                           | inst_eret             | inst_mtc0             | inst_addu | inst_sub             | inst_sltu | inst_multu | inst_bgez | inst_bgtz                         | inst_bgezal                          | inst_nor             | inst_or                        | inst_sra | inst_sllv             | inst_srav             | inst_mtlo | inst_lh | inst_sh | inst_lbu            | inst_jalr | inst_divu| inst_break); // 0

    // �Ƿ����ڴ�õ�������д�Ĵ���?
    assign id_mreg_o       = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu;
    
    // дHILO�Ĵ���ʹ���ź�
    assign id_whilo_o      = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_mult | inst_multu | inst_div | inst_divu | inst_mthi | inst_mtlo);
    
    // дͨ�üĴ���ʹ���ź�
    assign id_wreg_o       = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : jal ? `WRITE_ENABLE :
                             (inst_add | inst_subu | inst_and | inst_slt | inst_addu | inst_sub | inst_sltu | inst_or | inst_xor | inst_nor | inst_addiu | inst_ori | inst_sltiu | inst_lui | inst_addi | inst_slti | inst_andi | inst_xori | inst_mfhi | inst_mflo | inst_sll | inst_srl | inst_sra | inst_sllv | inst_srlv | inst_srav | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_mfc0 | inst_jalr);
    // ��ͨ�üĴ����Ѷ˿�1ʹ���ź�
    assign rreg1 = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_add | inst_subu | inst_and | inst_slt | inst_addu | inst_sub | inst_sltu | inst_or | inst_xor | inst_nor | inst_addiu | inst_ori | inst_sltiu | inst_lui | inst_addi | inst_slti | inst_andi | inst_xori | inst_mult | inst_multu | inst_div | inst_divu | inst_sllv | inst_srlv | inst_srav | inst_mthi | inst_mtlo | inst_lb | inst_lw | inst_lh | inst_lbu | inst_lhu | inst_sb | inst_sw | inst_sh | inst_jr | inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal | inst_jalr) & ~inst_lui;
    
    // ��ͨ�üĴ����Ѷ��˿�2ʹ���ź�
    assign rreg2 = (cpu_rst_n == `RST_ENABLE) ? 1'b0 : (inst_add | inst_subu | inst_and | inst_slt | inst_addu | inst_sub | inst_sltu | inst_or | inst_xor | inst_nor | inst_mult | inst_multu | inst_div | inst_divu | inst_sll | inst_srl | inst_sra | inst_sllv | inst_srlv | inst_srav | inst_sb | inst_sw | inst_sh | inst_beq | inst_bne | inst_mtc0);
    
    // ����ǰ�ƿ����ź�
    assign fwrd1[0] = (exe2id_wreg == `WRITE_ENABLE) & (exe2id_wa == rs);
    assign fwrd1[1] = (mem2id_wreg == `WRITE_ENABLE) & (mem2id_wa == rs);
    assign fwrd2[0] = (exe2id_wreg == `WRITE_ENABLE) & (exe2id_wa == rt);
    assign fwrd2[1] = (mem2id_wreg == `WRITE_ENABLE) & (mem2id_wa == rt);
    /*------------------------------------------------------------------------------*/

    // ��ͨ�üĴ����Ѷ˿�1�ĵ�ַΪrs�ֶΣ����˿�2�ĵ�ַΪrt�ֶ�
    assign ra1   = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD : rs;
    assign ra2   = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD : rt;
                                            
    // ��ô�д��Ŀ�ļĴ����ĵ�ַ��rt��rd��
    assign id_wa_o      = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD :
                          (jal) ? 5'b11111 :
                          (rtsel) ? rt : rd;

    // ���Դ������?1�����shift�ź���Ч����Դ������1Ϊ��λλ��������Ϊ�Ӷ�ͨ�üĴ����Ѷ˿�1��õ�����?
    assign id_src1_o = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD :
                       (inst_sll | inst_srl | inst_sra) ? sa :
                       (rreg1 == `READ_DISABLE) ? `ZERO_WORD :
                       (fwrd1[0] == 1'b1) ? exe2id_wd :
                       (fwrd1[1] == 1'b1) ? mem2id_wd : rd1;

    // ���Դ������?2�����immsel�ź���Ч����Դ������1Ϊ������������Ϊ�Ӷ�ͨ�üĴ����Ѷ˿�2��õ�����?
    assign id_src2_o = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD :
                       (immsel) ? imm_ext :
                       (rreg2 == `READ_DISABLE) ? `ZERO_WORD :
                       (fwrd2[0] == 1'b1) ? exe2id_wd :
                       (fwrd2[1] == 1'b1) ? mem2id_wd : rd2;
    
    assign id_din_o = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD :
                      (inst_sb | inst_sw | inst_sh) ? 
                      ((rreg2 == `READ_DISABLE) ? `ZERO_WORD :
                      (fwrd2[0] == 1'b1) ? exe2id_wd :
                      (fwrd2[1] == 1'b1) ? mem2id_wd : rd2) : `ZERO_WORD;
                      
                      
    assign id_retaddr_o = (cpu_rst_n == `RST_ENABLE) ? `ZERO_WORD : (id_pc_i + 8);
                      
    assign equ = inst_beq ? id_src1_o == id_src2_o :
                 inst_bne ? id_src1_o != id_src2_o :
                 inst_bgtz ? $signed(id_src1_o) > $signed(0) :
                 inst_blez ? $signed(id_src1_o) <= $signed(0) :
                 (inst_bgez | inst_bgezal) ? ~id_src1_o[31] :
                 (inst_bltz | inst_bltzal) ?  id_src1_o[31] : 1'b0;
    assign jtsel[1] = inst_jr | inst_jalr | ((inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal) & equ);
    assign jtsel[0] = inst_j | inst_jal | ((inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal) & equ);
    
    assign jump_addr_1 = {pc_next[31:28], instr_index, 2'b00};        //J, JAL
    assign jump_addr_2 = pc_next + { { 14 {imm[15]} }, imm, 2'b00};   //BEQ,BNE 
    assign jump_addr_3 = id_src1_o;                                   //JR,JALR
    
    assign stallreq_id = (cpu_rst_n == `RST_ENABLE) ? `NOSTOP :
                         (((exe2id_wreg == `WRITE_ENABLE && exe2id_wa == ra1 && rreg1 == `READ_ENABLE) ||
                         (exe2id_wreg == `WRITE_ENABLE && exe2id_wa == ra2 && rreg2 == `READ_ENABLE)) && (exe2id_mreg == `TRUE_V)) ? `STOP :
                         (((mem2id_wreg == `WRITE_ENABLE && mem2id_wa == ra1 && rreg1 == `READ_ENABLE) ||
                         (mem2id_wreg == `WRITE_ENABLE && mem2id_wa == ra2 && rreg2 == `READ_ENABLE)) && (mem2id_mreg == `TRUE_V)) ? `STOP : `NOSTOP;

    //�ж���һ��ָ���Ƿ����ӳٲ�ָ��                     
    assign next_delay_o = (cpu_rst_n == `RST_ENABLE) ? `FALSE_V : (inst_j | inst_jal | inst_jr | inst_jalr | inst_beq | inst_bne | inst_bgez | inst_bgtz | inst_blez | inst_bltz | inst_bgezal | inst_bltzal);
    
    //�жϵ�ǰ��������׶�ָ���Ƿ�����쳣����������Ӧ���쳣���ͱ���  
    assign id_exccode_o = (cpu_rst_n == `RST_ENABLE) ? `EXC_NONE :
                          (id_aluop_o == 8'h00) ? `EXC_RI :      //����δ����ָ��
                          (inst_syscall == `TRUE_V ) ? `EXC_SYS :
                          (inst_break == `TRUE_V) ? `EXC_BREAK :
                          (inst_eret == `TRUE_V ) ? `EXC_ERET : `EXC_NONE;
                          
    assign cp0_addr = (cpu_rst_n == `RST_ENABLE) ? `REG_NOP : rd;  //cp0�Ĵ������ʵ�ַ

endmodule
